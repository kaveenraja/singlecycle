module set(Of, Cf, Zf, Sf, Oper, out);
input Of, Cf, Zf, Sf;
input [3:0] Oper;
output out;

endmodule
